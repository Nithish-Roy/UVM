//interface.sv
interface seq_interface(input logic clk);

    logic        rst    ;
    logic        i_bit  ;
    logic        flag   ;

endinterface

