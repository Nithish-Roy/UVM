/***********************************************************************
************************UVM_PACKAGES_IMPORTING**************************
***********************************************************************/

`timescale 1ns/1ps

`include "uvm_macros.svh"

import uvm_pkg::*;

  /***********************************************************************
  ************************INCLUDING        FILES**************************
  ***********************************************************************/

	`include "interface.sv"
	`include "sequence_item.sv"
	`include "sequence.sv"
	`include "sequencer.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "agent.sv"
	`include "scoreboard.sv"
	`include "environment.sv"
	`include "test.sv"


  /***********************************************************************
  ************************TOP**************MODULE*************************
  ***********************************************************************/

module top;

  bit clk;
  
  alu_interface inf (.clk(clk));
  
  alu dut(
    .clock(inf.clk),
    .reset(inf.reset),
    .A(inf.A),
    .B(inf.B),
    .ALU_Sel(inf.select_line),
    .ALU_Out(inf.out),
    .CarryOut(inf.carry)
  );
  
  /***********************************************************************
  ****************************CLOCK GENERATION****************************
  ***********************************************************************/
  
  always #2 clk = !clk;
  
  initial begin
    
    $dumpfile("dump.vcd");
    
    $dumpvars();
    
  end
  
  
  /***********************************************************************
  ************************INTERFACE CONFIGURATION*************************
  ***********************************************************************/
  
  initial begin 
    
    uvm_config_db #(virtual alu_interface)::set(null,"*","vif", inf);
    
  end
  
  /***********************************************************************
  ********************************TEST RUN********************************
  ***********************************************************************/
  
  initial begin 
    
    run_test("alu_test");
    
  end
  
  /***********************************************************************
  ************************TERMINATE SIMULATION****************************
  ***********************************************************************/
  
  
  initial begin 
    
    #5000;
    
    $display("clock ended");
    
    $finish();
    
  end
  
endmodule
